library verilog;
use verylog.vl_types.all;
entity eyulingo_ios_dev is
    iter1(
        - [ ] 快速进入／退出 CartPageView 闪退问题
        - [ ] 点击购物车项目不能进入商品详情问题
        - [ ] 点击表头不能进入商店详情问题
        - [ ] 在短时间内（一分钟）没有进行购物车更新的情况下不要重复加载
        - [ ] 下拉更新，包括搜索页面以及购物车页面，以及将来的已购商品页面
        - [ ] CI/CD
    );
end eyulingo_ios_dev;